`default_nettype none

// Fetches the background tiles from memory.
// https://gbdev.io/pandocs/pixel_fifo.html
// https://hacktix.github.io/GBEDG/ppu/#background-pixel-fetching
module BackgroundFetcher #(
    parameter X_MAX = 160,
    parameter TOTAL_SCANLINES = 154
) (
    // Standard clock and reset signals.
    input wire clk_in,
    input wire rst_in,

    // The T-cycle clock.
    input wire tclk_in,

    // Access to the internal X position counter.
    input wire [$clog2(X_MAX)-1:0] X_in,
    // Access to the internal Y position counter.
    input wire [$clog2(TOTAL_SCANLINES)-1:0] Y_in,

    // Access to the SCY and SCX registers.
    input wire [7:0] SCY_in,
    input wire [7:0] SCX_in,
    // Flag to determine which background map to use for the background.
    input wire background_map_in,

    // Access to the WY and WX registers.
    input wire [7:0] WY_in,
    input wire [7:0] WX_in,
    // Determines if the WY condition is met.
    // https://gbdev.io/pandocs/Scrolling.html#ff4aff4b--wy-wx-window-y-position-x-position-plus-7
    input wire WY_cond_in,
    // Flag to determine which background map to use for the window.
    input wire window_map_in,
    // Flag to determine if the window is enabled.
    input wire window_ena_in,

    // Determines which addressing scheme to use for accessing background tiles.
    input wire addressing_mode_in,

    // Wire requesting a tile row from memory.
    output logic [15:0] addr_out,
    // Valid request to fetch data from memory.
    output logic addr_valid_out,
    // Data fetched from memory.
    input wire [7:0] data_in,
    // Whether the data fetched is valid.
    input wire data_valid_in,

    // Wire to tell the fetcher has completed a pixel push to LCD.
    output logic advance_X_out    
);
    // Defines the 4 states that takes 2 T-cycles each.
    typedef enum logic[1:0] {
        FetchTileNum = 0, 
        FetchTileDataLow = 1, 
        FetchTileDataHigh = 2, 
        Push2FIFO = 3
    } FetcherState;
    FetcherState state;
    // Determines whether or not we are waiting a T-cycle to advance the state.
    logic stall;
    // Counts the number of elapsed T-cycles.
    evt_counter #(
        .MAX_COUNT(2)
    ) evt_counter (
        .clk_in(tclk_in),
        .rst_in(rst_in),
        .evt_in(tclk_in),
        .count_out(stall)
    );

    // The state evolution of the fetcher.
    always_ff @(posedge tclk_in && stall) begin
        if (rst_in) begin
            state <= FetchTileNum;
            addr_out <= 16'h0;
            addr_valid_out <= 1'b0;
            advance_X_out <= 1'b0;
        end else begin
            case (state)
                FetchTileNum: begin
                    if (X_in == $clog2(X_MAX)'(X_MAX-1)) begin
                        state <= FetchTileDataLow;
                    end
                end
                FetchTileDataLow: begin
                    state <= FetchTileDataHigh;
                end
                FetchTileDataHigh: begin
                    state <= Push2FIFO;
                end
                Push2FIFO: begin
                    state <= FetchTileNum;
                end
            endcase
        end
    end

    // Tracks the X position of the fetcher within the tile.
    logic [$clog2(31)-1:0] fetcher_x;
    logic x_progress;
    evt_counter #(
        .MAX_COUNT(32)
    ) tile_x_counter (
        .clk_in(tclk_in),
        .rst_in(rst_in),
        .evt_in(x_progress),
        .count_out(fetcher_x)
    );
    // Tracks the Y position of the fetcher within the tile.
    logic [$clog2(255)-1:0] fetcher_y;
    logic y_progress;
    evt_counter #(
        .MAX_COUNT(256)
    ) tile_y_counter (
        .clk_in(tclk_in),
        .rst_in(rst_in),
        .evt_in(y_progress),
        .count_out(fetcher_y)
    );

    // Combinational logic determining if we are inside of a window.
    logic inside_window;
    assign inside_window = (X_in + 7) >= WX_in && window_ena_in && WY_cond_in;
    // Tracks the window tile X position.
    logic [$clog2(31)-1:0] window_tile_x;
    evt_counter #(
        .MAX_COUNT(32)
    ) window_x_counter (
        .clk_in(tclk_in),
        .rst_in(rst_in),
        .evt_in(x_progress && inside_window),
        .count_out(window_tile_x)
    );
    // Tracks the window Y position.
    logic [$clog2(255) - 1:0] window_y;
    assign window_y = (WY_in - Y_in) & 8'hFF;

    // Determines the base tile address to fetch from.
    logic [15:0] base_addr;
    always_comb begin
        // Determines the base address to fetch from.
        if (background_map_in && !inside_window) begin
            base_addr = 16'h9C00;
        end else if (window_map_in && inside_window) begin
            base_addr = 16'h9C00;
        end else begin
            base_addr = 16'h9800;
        end
    end
    // Determines the offset from the base address to fetch the tile number from.
    logic [9:0] tile_offset;
    // Fetches the tile number to request.
    logic [7:0] tile_num;
    assign tile_offset = (SCY_in + Y_in) & 8'hFF;
    always_ff @(posedge tclk_in) begin
        if (rst_in) begin
            tile_num <= 8'h0;
        end else begin
            if (state == FetchTileNum) begin
                // First cycle make address request.
                if (!stall) begin
                    if (tclk_in) begin
                        addr_out <= base_addr + tile_offset;
                        addr_valid_out <= 1'b1;
                    end
                // Second cycle save the tile number.
                end else begin
                    if (data_valid_in) begin
                        tile_num <= data_in;
                    end
                    addr_valid_out <= 1'b0;
                end
            end
        end
    end

    // Tracks the address base of the tile.
    logic [15:0] tile_addr;
    always_comb begin
        tile_addr = addressing_mode_in ? 
            (16'h8000 + (12'(tile_num) << 4)) : 
            (16'h9000 + (12'($signed(tile_num)) << 4));
    end
    // Tracks the low byte of the tile data.
    logic [7:0] tile_data_low;
    always_ff @(posedge tclk_in) begin
        if (rst_in) begin
            tile_data_low <= 8'h0;
        end else begin
            if (state == FetchTileDataLow) begin
                // First cycle make address request.
                if (!stall) begin
                    addr_out <= tile_addr;
                    addr_valid_out <= 1'b1;
                end else begin
                    if (data_valid_in) begin
                        tile_data_low <= data_in;
                    end
                    addr_valid_out <= 1'b0;
                end
            end
        end
    end

    // Push2FIFO state logic.
    always_ff @(posedge tclk_in) begin
        if (rst_in) begin
            advance_X_out <= 1'b0;
        end else begin
            if (state == Push2FIFO && !stall) begin
                advance_X_out <= 1'b1;
            end else begin
                advance_X_out <= 1'b0;
            end
        end
    end
endmodule

`default_nettype wire